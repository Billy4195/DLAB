`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:03:13 12/26/2015 
// Design Name: 
// Module Name:    final_pro 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module final_pro(
    input  clk,
    input  reset,
    input start,
	 input ROT_A,
	 input ROT_B,
    //input  [1:0] button,

    // VGA specific I/O ports
	 output reg [7:0] led,
    output HSYNC,
    output VSYNC,
    output VGA_RED,
    output VGA_GREEN,
    output VGA_BLUE
	);
	
	// general VGA control signals
wire video_on;      // when video_on is 0, the VGA controller is sending
                    // synchronization signals to the display device.

wire pixel_tick;    // when pixel tick is 1, we must update the RGB value
                    // based for the new coordinate (pixel_x, pixel_y)

wire [9:0] pixel_x; // x coordinate of the next pixel (between 0 ~ 639) 
wire [9:0] pixel_y; // y coordinate of the next pixel (between 0 ~ 479)

reg [2:0] rgb_reg;  // RGB value for the current pixel
reg [2:0] rgb_next; // RGB value for the next pixel

// Application-specific VGA signals
wire [2:0] current_rgb; // RGB values for the frame display application.
                        // In this demo, the value is generated by
                        // a video pattern generator:
                        //      video_pattern(id, x, y, current_rgb),
                        // where the input is the current scan coordinate (x, y),
                        // and the output is the RGB value of the video pattern
                        // 'id' at pixel (x, y).
reg start_b;
								
reg [9:0]gp_pos_x;
reg [9:0]gp_pos_y;

reg [9:0]tp_pos_x;
reg [9:0]tp_pos_y;
reg tp_show;
reg [3:0]tp_cnt;
reg [1:0]tp_id;

reg fb_show;
reg [2:0]score;

wire [2:0] rgb_gp;
wire [2:0] rgb_stbd;
wire [2:0] rgb_tp;
wire [2:0] rgb_fb;

reg [3:0]score_0;
reg [3:0]score_1;
reg [3:0]score_2;
reg [3:0]score_3;

reg led_valid;
reg catch;

localparam init_s = 3'b000 , set_s = 3'b001,fall_s = 3'b010 , dsap_s = 3'b011 , over_s = 3'b100;

reg [2:0]S_cur,S_next;

//reg [25:0] cnt;
reg [19:0] cnt;
reg [25:0]rand;

// Declare system variables
//wire [1:0]  btn_level, btn_pressed;
//reg  [1:0]  prev_btn_level;	

wire stbd_valid;
wire gp_valid;
wire tp_valid;
wire fb_valid;		

//debounce btn_db0(
//  .clk(clk),
//  .btn_input(button[0]),
//  .btn_output(btn_level[0])
//  );
//
//debounce btn_db1(
//  .clk(clk),
//  .btn_input(button[1]),
//  .btn_output(btn_level[1])
//  );

// instiantiate a VGA sync signal generator

initial begin
	gp_pos_x = 319;
	gp_pos_y = 463;
	tp_pos_x = 319;
	tp_pos_y = 10;
   start_b = 0;
   tp_show = 0;
end
vga_sync vs0(
  .clk(clk), .reset(reset), .oHS(HSYNC), .oVS(VSYNC),
  .visible(video_on), .p_tick(pixel_tick),
  .pixel_x(pixel_x), .pixel_y(pixel_y)
  );
  
GP gp(
	.clk(clk),
	.midx(gp_pos_x),
	.midy(gp_pos_y),
	.x(pixel_x),
	.y(pixel_y),
	.rgb(rgb_gp),
	.gp_valid(gp_valid)
    );

TP tp(
	.clk(clk),
	.show(tp_show),
	.id(tp_id),
	.midx(tp_pos_x),
	.midy(tp_pos_y),
	.x(pixel_x),
	.y(pixel_y),
	.rgb(rgb_tp),
	.tp_valid(tp_valid)
    );
	 
status_board sta_bd(
	.x(pixel_x),
	.y(pixel_y),
	.id(tp_cnt),
	.rgb(rgb_stbd),
	.stbd_valid(stbd_valid)
    );
Rotation_direction rd(
    .CLK(clk),
    .ROT_A(ROT_A),
    .ROT_B(ROT_B),
    .rotary_event(ro_event),
    .rotary_right(ro_dir)
    );
final_board fb(
    .clk(clk),
    .show(fb_show),
    .score_0(score_0),
    .score_1(score_1),
    .score_2(score_2),
    .score_3(score_3),
	 .x(pixel_x),
	 .y(pixel_y),
	 .rgb(rgb_fb),
	 .fb_valid(fb_valid)
    );

// Button click controller
//always @(posedge clk) begin
//  if (reset)
//    prev_btn_level <= 2'b11;
//  else
//    prev_btn_level <= btn_level;
//end
//
//assign btn_pressed = (btn_level & ~prev_btn_level);

// VGA color pixel generator
assign {VGA_RED, VGA_GREEN, VGA_BLUE} = rgb_reg;

//init 
always@(posedge clk)begin
   if(start)
      start_b <= 1;
   else 
      start_b <= 0;
end
always@(posedge clk)begin
   if(start_b)
      S_cur <= init_s;
   else begin
      S_cur <= S_next;
   end
end

//state control
always@(posedge clk)begin
   case(S_cur)
   init_s:
      S_next <= set_s;
   set_s:
      S_next <= fall_s;
   fall_s:
      if(catch || tp_pos_y >= 470)
         S_next <= dsap_s;
      else
         S_next <= fall_s;
   dsap_s:
      if(tp_cnt == 0)
         S_next <= over_s;
      else 
         S_next <= set_s;
   over_s:
      S_next <= over_s;


   endcase

end

always @(posedge clk) begin
  if (pixel_tick)
    rgb_reg <= rgb_next;
  else
    rgb_reg <= rgb_reg;
end

always @(*) begin
  if (~video_on)
    rgb_next = 3'b000; // synchronization period, no need to set RGB values
  else
    rgb_next = current_rgb; // RGB value at (pixel_x, pixel_y)
end
	
assign current_rgb = stbd_valid ? rgb_stbd: gp_valid ? rgb_gp : tp_valid ? rgb_tp : fb_valid ? rgb_fb : 111;
//assign rgb_gp = 3'b000;
//assign rgb_stbd = 3'b000;

//GP controller
always@(posedge clk)begin
	if(S_cur == init_s)begin
		gp_pos_x <= 319;
		gp_pos_y <= 463;
	end
	else if(ro_event)begin
		if(ro_dir)begin			//right
			if(gp_pos_x <= 619)
				gp_pos_x <= gp_pos_x + 20 ;
			else
				gp_pos_x <= 639;
		end
		else begin					//left
			if(gp_pos_x >= 20)
				gp_pos_x <= gp_pos_x - 20;
			else
				gp_pos_x <= 0;
		end
	end 
end

//TP controller
always@(posedge clk)begin
	if(S_cur == init_s || S_cur == set_s)begin
		tp_pos_x = 0 + 30 *(rand % 16);
		tp_pos_y = 10 + 10 * (rand % 8);
		tp_show <= 1;
		tp_id = rand % 4;
	end
	else if(S_cur == fall_s)
      if(cnt == 1000000)begin
         if(tp_pos_y < 479)begin
            tp_pos_y = tp_pos_y + 4;
            tp_show <= 1;
         end
         else
            tp_show <= 0;
      end
 
end

//TP conunter
always@(posedge clk)begin
	if(S_cur == init_s)
		tp_cnt <= 10;
   else if(S_cur == set_s && S_next == fall_s)
      tp_cnt <= tp_cnt -1;

end

//cnt counter
always@(posedge clk)begin
//	if(S_cur == init_s)
//		cnt <= 0;
//	else 
   if(cnt < 1000000) //1 million
		cnt <= cnt + 1;
	else
		cnt <=0;

end


always@(*)begin
   if(rand < 1500000)
      rand <= rand + 1;
   else 
      rand <= 0;
end

//collision handler
always@(posedge clk)begin
	if(S_cur == init_s)begin
//		led <= 8'd0;
//		led_valid <= 1;
      catch <=0;
	end
	else if(S_cur == fall_s)begin
				if(tp_pos_x <= gp_pos_x+10 && tp_pos_x >= gp_pos_x-10 && tp_pos_y <= gp_pos_y+10 && tp_pos_y >= gp_pos_y-10)begin
//					led <= led + 1;
//					led_valid <= 0;
               catch <= 1;
				end		
			end
         else if(S_cur == dsap_s)
            catch <=0;
end

//led 
always@(posedge clk)begin
   if(S_cur == init_s)begin
      led <= 0;
      score_0 <= 0;
      score_1 <= 0;
      score_2 <= 0;
      score_3 <= 0;
   end
   else if(catch && led_valid)
      led <= led + 1;
      case(tp_id)
      0:score_0 <= score_0+1;
      1:score_1 <= score_1+1;
      2:score_2 <= score_2+1;
      3:score_3 <= score_3+1;
      endcase
//   else
//      led <= tp_cnt;
end
always@(posedge clk)begin
   if(S_cur == set_s)begin
      led_valid <= 1;
   end
   else if(catch)
      led_valid <= 0;
end
//final board 
always@(posedge clk)begin
   if(S_cur == over_s)begin
      fb_show <= 1;
   end
   else
      fb_show <= 0;
end

endmodule
